module AND_bitwise(data_operandA, data_operandB, result);

   input [31:0] data_operandA, data_operandB;

   output [31:0] result;

	and and_g0(result[0], data_operandA[0], data_operandB[0]);
	and and_g1(result[1], data_operandA[1], data_operandB[1]);
	and and_g2(result[2], data_operandA[2], data_operandB[2]);
	and and_g3(result[3], data_operandA[3], data_operandB[3]);
	and and_g4(result[4], data_operandA[4], data_operandB[4]);
	and and_g5(result[5], data_operandA[5], data_operandB[5]);
	and and_g6(result[6], data_operandA[6], data_operandB[6]);
	and and_g7(result[7], data_operandA[7], data_operandB[7]);
	and and_g8(result[8], data_operandA[8], data_operandB[8]);
	and and_g9(result[9], data_operandA[9], data_operandB[9]);	
	and and_g10(result[10], data_operandA[10], data_operandB[10]);
	and and_g11(result[11], data_operandA[11], data_operandB[11]);
	and and_g12(result[12], data_operandA[12], data_operandB[12]);
	and and_g13(result[13], data_operandA[13], data_operandB[13]);
	and and_g14(result[14], data_operandA[14], data_operandB[14]);
	and and_g15(result[15], data_operandA[15], data_operandB[15]);
	and and_g16(result[16], data_operandA[16], data_operandB[16]);
	and and_g17(result[17], data_operandA[17], data_operandB[17]);
	and and_g18(result[18], data_operandA[18], data_operandB[18]);
	and and_g19(result[19], data_operandA[19], data_operandB[19]);
	and and_g20(result[20], data_operandA[20], data_operandB[20]);
	and and_g21(result[21], data_operandA[21], data_operandB[21]);
	and and_g22(result[22], data_operandA[22], data_operandB[22]);
	and and_g23(result[23], data_operandA[23], data_operandB[23]);
	and and_g24(result[24], data_operandA[24], data_operandB[24]);
	and and_g25(result[25], data_operandA[25], data_operandB[25]);
	and and_g26(result[26], data_operandA[26], data_operandB[26]);
	and and_g27(result[27], data_operandA[27], data_operandB[27]);
	and and_g28(result[28], data_operandA[28], data_operandB[28]);
	and and_g29(result[29], data_operandA[29], data_operandB[29]);
	and and_g30(result[30], data_operandA[30], data_operandB[30]);
	and and_g31(result[31], data_operandA[31], data_operandB[31]);


endmodule
